`timescale 1ns / 1ps
/**
 * Copyright: Steven van der Schoot
 */
module stress(
    input  [7:0] hartvolume,
    input  [7:0] huilvolume,
    output [7:0] stress
    );
	
	
	
endmodule
