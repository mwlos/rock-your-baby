module hoogLaag()

endmodule
