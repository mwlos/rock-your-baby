module holdReset(
	input clk,
	input resetSignal,
	input stopHold,
	output reset);
	
	
	
endmodule
