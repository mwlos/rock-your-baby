module huilVolume(
	input clk,
	input slowClk,
	input reset,
	input [7:0] DSPinvoer,
	input DSPready,
	output reg [7:0] huilVolume);
	
		
	
endmodule
